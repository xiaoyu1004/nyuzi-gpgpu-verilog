`ifndef DEFINES_VH
`define DEFINES_VH

// `define VENDOR_XILINX

`endif