`include "defines.vh"

module ifetch_tag_stage(
    input                           clk             ,
    input                           rst_n           ,
);
endmodule