`ifndef DEFINES_VH
`define DEFINES_VH

`define SIMULATION
`define ENABLE_SV_ASSERTION

`endif