`ifndef CONFIG_VH
`define CONFIG_VH

parameter NUM_VECTOR_LANES  = 16;

parameter L1_CACHE_NUM_WAYS   = 4;
parameter L1_CACHE_NUM_SETS   = 16;


`endif